module mux16bit221(
    input [15:0] A,
    input [15:0] B,
    input sel,
    output reg [15:0] out
);

always @(*) begin
    case (sel)
        0: out = A;
        1: out = B;
        default: out = A;
    endcase
end

endmodule