`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:20:47 11/26/2023 
// Design Name: 
// Module Name:    adder16bit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module adder16bit(
    input [15:0] A,
    input [15:0] B,
    output reg [15:0] S
    );
always @* begin
    S = A + B;
end

endmodule
